PK   �DV)�U�#  �\    cirkitFile.json�O��F�ſ��s�FGeU�n;�q�3v�7<I� �bL��e�-{��[	v�I�:_����-����D�P����տv��z��_���f{�zE���]�k?�ǯ��Շ�m��V����V�>������uu�l�>պ����"Y��$�%u�MR���Z���u_�ʬ^�~{�r+���RSY1�T�TN� U0�3HL���
���RS�b���
1�T�T��A�j��P�%�T�k%ɋ�X"P�˥X"P��X"P�K�X"Pȋ�X"P�˦X"P��X"P�K�X"���S,(�S,( My���)���)���)���)���)���)���)��P^;��B^;��B^;��`����k�X"P�k�X"P�k�X"P�k�X"P�k�X"P�k�X�T^^;��B^;��B^;��B^;��p�S^;��v�%��v�%��v�%��v�%��v�%L��k�X"P�k�X"P�k�X"P�k�X"P�k�X"P n�kg*��b�@!��b�@!��b�@!��b	Se��)���)���I|�~�vɮ��̞�P}��Ի�����R��E(GX:�ҙ �ac�#,��,6v;(a�L就s��A�K<6v;(a���;(a����;(a�L�cc�cc�#,��
l�
l�t��3U��]�����t<+<8;,��x>#8~hw��`A`�A`���#0�!��2�|��ٯ�������|<o?������g��vX>��\ip����G`>����y`��������,��xf=�3�`���k�|Oj������v_e�<oK�	G��m�֦�);�LY�����z�u���B�9�O�ښ�Y'y���wm��}�'mf|�e��uV�4���*�+`�c#W���[i���)�j8=H�#C��CF{�ي�N{�ٲ`���#0/Q�l��|t����j)=T#��-�`�5�$��ς-���|��?������ ����-���|�t?�O����]��6[X>��rQp����3���Ɂo19���������v=1߹�-9�]o�$�|���̓�ͳ��e���m	��x]28�`��}���(O���|MRfe�ؾ����+3#�G�Ƌ����,��{�O)5�l��0a���k���&,��{�%Qa�z���`���#0�: �쵰|��&�������|�^?������c��^8�^9�Z�<�ka����H��&,����
8~`׃�3|/:�ҡ#��x�������ހ�v=X>�q�l�R�u����;���.X>�q�$p����G`>���غ`���}���[,����8~���`뒂�K
�.X>�q3p����G`>���`��ǝ����,����6~�`��������,���� 8~`���|G�z�ue�&�/�ܺ���]R�]ӧ.�����p�q�ȅ���;.�}��v���f�ww�]��������}[�>n��p�q�ԥi#M;a�EϠ[��0��-�_�{ѳ֖�/̾��fK��_�L���K�0��'p-�_��S���/̿�ISK��_�t��'.a�EOTZx�뙏�7���v�|ޗ �i���Gsv��g�Y&��~� �ײ@���(�0��w�(�T�yK=e�d��Tr������3���E
C���u��>���V�0+�gN��ds~��+��Y��PdQ���P�et���灥�o���f�[���$����G[��VW/"�А�"���C2<�����0D !Ã*H��8C2<\�����0D !�AH��AP��Um\ن�m�n��.6��`��`��d��� &X�&XG)���-�	V�	V�QJf��b��q��(%3\1��߸8��[XG)��F �	V�-�����p����V�QJf��b��q��(%3� �qXw�:�R�Q0&ܕܥXw�:�R�vA0&Xw�:�R�30&Xw�:�R�n&0&X��:�R��0&X��:�R�0&�5q�EqX��:�R���0&X��:�R��0&X��:�R�5ϰ[?�:���8J���`u<��q��!�1��n�no��x
��(%^?c���V�QJ���������x=�	V�3X�RZ>mi�L�:,�B��
+���j�|�
��+���j���
��+���j�n�
��+��ߥ�q3L4XI�5��T�:nR���+���1�J\��K0�`%VS�ۙ�U�q�`%VS�ۜ�U�q�`%VS�۟�U�q�`%V��ct�
-����f��*�.%ۥ�H�x���R�%Z�k�[��BK:�<g^'�:L��thy�Nlu\�
-������81Zҡ�:��qc*��C�kJtb���ThI������VǕ�В-��ѹ����ThI�6�[d��+����/S��;`�b�tGL閘�/��@�VǗ��E�"c;Hlu|�Z�,2�:����2Zҡ5'����e*�qϴA6O�A���&���3�hYd���2���ThI��׺��VǗ�В-��ՙ����ThI�����VǗ�В-��։��/S�%Z^�[�يJ�u|�ӹ_�t|�
-�К����,2�1�|4N:�&ꏫ ��mL����2�s�l�][_v�V�y��/s:�L��th������e*��c@y�u|���e*��C˽Dtb���ThI��{���VǗ�В-�vщ��/S�%Z�Q�[��dJK�t|���e^Ǘ�В-�҉��/S�%Zs�&dlu|�
m�$*��VǗy_�BK:�܋J'�:�L��th���JlS_�BK:��L'�:�L��th�ǙNlu|�
-��r�6����2Zҡ�s:���e*��C˽�tb���C�͇�/Ku|Y���ThI��{��VǗ�В-�dԉ��/S�%Z�-�[_�BK:��#S%���/S�%Z���[_�BK:�ܳT'�:�L����=ؼwYWvi��"���>)m�%u�5}�R�����0/T��M�Pe���B��>�U&:o/T�蕽Pe���B��~�U&:H/T����4�@ɋ�ީ��.����ԣU��`2x��Ke09<��Х2�,�z�RP�d��S*��`�x�Y�Ke0Y<��ť2�,�z��ҳ.&���x$���ta��QвM�[�&��3e�n�vƨf�
����P��5G���4G�p8�1Y.P�|4�Q�x��B��]>�樔�è������&O�η���<��<KZ[�o��i�
�B��ڬ&Gy��]���M�2+����-�u]ܶ��Y*t��~mM٬����Ļ6��M����Y�Y�����R���#�σL��Vw�z߭^}z�]�������~W��-�H���A�@Bf�>�$d�"!	��!	���!	��D!	��!	��!	��d!	�ÉS"qUW�au�`��dWm0L��M��R2��I&X�&XG)�Õ.���������	V�-������� �	7���au���8J�.�b�`u���8J�.�b�`u���8J�.c�`u���8J�.ic�8��;XG)q3(�J
�R
��;XG)q���;XG)q���;XG)qS��{XG)q��{XG)q��8�8��{XG)��x��{XG)�bl��{XG)��_حXOau�ċMaL�:���8J�7pw7q�7au<��q�/B�1��x
��(%^�c���V�QJ�������O)-_0-�B�ֵ TI��TXM-�B���J*���b�U�q�`%VSE�1Ъ��j��
k�]*q��b@"��J*�a�ר'$����(*q��a@"��J*����a�U�q�`%VSE�0Ъ��j��
���&hU`\5XI����ǥBK:�<�Y'�J�K�v��.�1^��ThI�����V�}�В-ϙ׉��S�%Z���[�BK:���A'�:NL��thy-�Nluܘ
-������82Zҡ�1:��qe*��C�k|tn,��2Zҡ�J:���e*��C�k�tb�tGL閘�/�:����2Zҡ�5p:���e*��C�k�tb���ThI���$��VǗ�В-��ԉ��/S�%Z^#�[_�BK:���U'�:�L��thyͮ��$_�BK:���X'�:�L��thy�Nlu|�
-���Zp��*�VT����˜�/s:�L��thym�Nlu|�
-��r�����2Zҡ�^	:���e*��C�=tb���ThI��{W��VǗ�В-��P����e*��C˽Dtb���ThI��{���VǗ�В-�vщ��/S�%Z�Q�[��dJK�t|���e^Ǘ�В-�҉��/S�%Z�}�[_�BK:���I'�:�L��th��Nlu|�
-��rO-�ئ:�L��th�7�Nlu|�
-��r�3����2Zҡ�^m:���e*��C�=�tb���ThI��{���V�ˇR�_����TǗ�В-�2ԉ��/S�%Z�ɨ[_�BK:��[R'�:�L��th�G�Jl3_�BK:���S'�:�L��th�g�Nlu|�
-ͣ=z*xﲮ����EP]w}RھK�k�ԥ>_7S�a^�2ћv��D7م*}��Lt�^�2�+{��Dw�*���Lt�^�2��yiց���S}]*��ߩG�.��d��L��`rx�1�Ke0Y<�0Υ2���⩧T.��d�Գ ��`�xꉋKe0Y<�\åg]LO==�Hf��m��~���e��6ML�Yg�r�4�Q���j����i����i���i���i���ci���Ci���#iV�]L^rֻ��I��6�Y�'u�gIkˢ�M�7M���r��6��Q�ty�'>|����:�}oKk]W�}�e��E�ԯ�)�u�y�x���ɓ63>�2��:��2K�r\>_������ۛ�ڴ��^����f��Un�u�V��j�k�����ׂ(�<�x��۫��!����	�|���Л�ʼCNRߥA]v��<'�0��CgcM��,�KL��ѱ7i��X!���2s !C!
I���XJ�!4n������h׽��NG�m{���:@��E���9�ɉ�g�3D����}�s&$�S߳!�C΀�C���/(]�@CN�oȉ���q�}ȉ��9|,�/r�����ջ�~s������[����m�~�j���7��է�w��H��Lu�˟C*�8\\R�%�pAHH!�0õf!�X�ת�b	3\�R�%�p�\H!�0õv!�X���b	3\�R�%��^��l!�'�|�'
�\�&qH9 5� ET�a�H��:J�B*�0��,R@-%@1�k��T)��Z@=�k��d)b<����S��9�G�r ��S��9̈�r ��S��9�ɒr ��S��9�
�ZI@=u�z*��� ��GX|@=u�z*��޵ @=u�z*���� @=u�z*��^� @=��z*��� @=��z*��ހ �5S�ES@=��z*���l @=��z*��_ @=��z*��~R����z��\��8 �4�S���p �B!nC�i
��r�A� ��PO���������5�g�PO3@=�5�O��h���Dz�#0���^8=H��|�3U������|��z�� ����/�p��F����#0__��5~_,���8 ��a���b��g��7 N?,��L����A��#0���8=H��|��y��4ځ�		M�s,�1���A�BB;0!�	yn+:�h7&$4!��E��H���&�9���]	��Є<C�3���r�c�v'`BB�<tt�LHhB�C��!ڥ�		M������>LHh�xE���9�#Z~��	)ڶ�	�F
QHE�BN�1!��PA��q'�(�NR���}#�!E�����q����}>B{0!�	�I�L�L�K��Dic��P����)���@AL���E; 0!�	y�:�h&$4!��CO5A; 0!�	y�!:�h�&$4!��D��q���&�U�����'��M�Cߩqh&$4����B11�GZQ�IB��O1T҈pRi_d�}���3��,)��Ą��H���8���М����mj��q'�(-�,�q<��		M� �1D{0!�	�{:�h�&$4!w^@��q���&������Ƞ=�G{��8`BBr�tѦLHhBs��L�.L?�$.���]�G�0!�	��:�h&$4!7��0E�0!�	��:�h�&$4!7	B�m[���&�G��m��Єܜ	C�m��K�c_�_ۏ�-)ڶ�h�&$4!7�B�m[���&�fd��}
��Є�HC�O�����c��}
��Є��C�O����c��)`B�Dx����e]٥������}��i���K}�n��*.�?j��p�����������.�?j��p��Q��������.�?j(�4�	(���YpK�9?}m��4��-��a�����L���T@\��?�j��4�N-�fb�����L�����&���1F�����Ǔ_�ϵP��b���s����q�玑y��~��B����ԅr�>�#��Rƥ�hb=s^����7y�w�M|V�I��Y�ڲh}��M�W�����rg���Ԣ6��Q�ty�'>|ɤ��:�}oKk]Wf��D�fɝ���]��֔�:ɋ�L�k�\��I��e��~����rg�r������Փ̦���*��i5��^�^q��G�4�ߖ+!`�ՙ����;���ěoK�1��ěoO������6�ay�{X���������=�No���8z�e��I���;��Ó�����a�<M��]bҾ�:O����d�6]�ٮ(�.��6����_����\�W�A>������]�t$��.�]���	�|����tn*v�d��xi�F�}%��.���At>XL�M��<Q�."�[�t��N���^�+$t�etqӞ���䝴k]���S�����_:7����q˒����m_��Mw�'����ƿw�o88�w��-�߲o��-����o�����4~+{x+�����㷊�������2z��Aq8�K8����Mu�,��m��n6w{N�Y?Y�*[����\�~ReMz�ɪ��q�G~�㻿��:|ا�w��n�������?N����ns˧���=��߽Z�Z����}P���v�W�ow���6�^���]޼�v?o�6�M��]�_��]����5��𾾽����~��8��d��on� ��j�f�ن8�N��.���*5�:O��kCd����Eۤ޸$�M�{�Nj�DѸ�J�����Ѿ�]��吮V��&�t�l����n^]ov����|�P�_�c�+_�o�ν���4�����O�M�O�QN�٩7�?��f����J����������G)blv�9٬��̧�6�����J3�+�&�����7\6�F:�����9�Ff҉7��g���f�����'�ɦs�E��v8�������o7۟��ݡ�5]�p;S�O���M���yam�<{�*�s>όˆ���XӅH��IҴ쓼E��އ3�w�7�񮉊؜�$�"�n?�F5̗�#�t�'4N�3[eٵ�e���㭊ö�|�	��6-3�o�l�<�ě9�Ct���vTPȪ����<���?�%(���c���#6�3�5���/�h�d��4_�V�ʺ�?��3��:#w(�g�Y宋4-J{x�m��uʰY�_ې�!��p�gƖ��E���|H�%�!E>\��Çm���7�o��m�y��>�#����$�P���<KS�E��xl]i��Mʴ���IYtu�^��m�v&:g]a�a�8>��塎>�ݚ봤��_!��������/2_>��UQҵ'�J*�SV�m��ƵI�0X��$�]�BNyZwy7FY1�2�H\`M��|S=�#�*mC��
y��_�
��H��|��f���C8]_��snB2�W�^��S����s������<Y��yєIY��~m�p�ѷ�8f�#�����w�����a�S���0�	y���r#��}�x��y������o��o��s��w�߿��_��)ʃǫ.G��/s�������g���Z�7��>Z�7�l��~����N������e���m���l��	f���w�S?�y�?��Çz}���}��V_>����U��O�QN��S����O���Ϊ~y��\T�T:B�v{��7�>>�wzS�cHD�̧&�����8jfa��NJ�O���&�+ˤ��'�+\�Q_���A':�gݳ�|_:*����p4��Zǣ{	Z7]�I҂��`(�:��M��
a�0�_9���.\�Z��aP^�m���'�|w�^���?�f�����y�}�G��_8��&ԍ�OoV�ެ���w���՛P)�]8�n�o��^|Cr�n�3R���������5��U��v�W�7�z��͊/b����o�4��;~��k��a��e�[���zÚ�f]��e�=���Yy�#�7z����sH���1Ç!��`����8y<y��J�'7�~��*/��|V,+)�n�c�"}iI�ϊ̊3��b0�O?df�� ��<s�ܟM�Q=�6��'dL�#3繓��)�D�p�y�0/��X���yv|���;�=��'�ڪ��n�z�|��8�������+��3�ܭN.j~����gj�n8�λ��-��O�X�e���Ã���9�p���[f�7��k�NM��q�V`��]�:O�5�˭�ӟ�զY[�sRg�VVaH7oN0��)r�l+,���.M0:I
��=�e�7ʢ�8�H����f_+s�g�h�"8s�g����y�=*Y�|�ԟM�q�ě}�ܱ��q��c�sW�;�7+FYA'q�Vi6��ěrg�\_l��sg+2w��`H4��jH�4��N~p��Ƴ.��mv�&O�cO�l�v�����f_+	<���H������8��!����&Zv����sY��=*�'�k�v���Q>F�}-�XB�hn?8K�a<��B����q�٩�4+�"l���_�=M�y[M\�x�C"���������}���7��(������w�������������wo�e����PK
   �DV)�U�#  �\                  cirkitFile.jsonPK      =   $    